module Sign32Bit(out,in);
    output [31:0] out;
    input [31:0] in;
    wire [31:0] S32Bcout;
    not n0(out[0],in[0]);
	not n1(out[1],in[1]);
	not n2(out[2],in[2]);
	not n3(out[3],in[3]);
	not n4(out[4],in[4]);
	not n5(out[5],in[5]);
	not n6(out[6],in[6]);
	not n7(out[7],in[7]);
	not n8(out[8],in[8]);
	not n9(out[9],in[9]);
	not n10(out[10],in[10]);
	not n11(out[11],in[11]);
	not n12(out[12],in[12]);
	not n13(out[13],in[13]);
	not n14(out[14],in[14]);
	not n15(out[15],in[15]);
	not n16(out[16],in[16]);
	not n17(out[17],in[17]);
	not n18(out[18],in[18]);
	not n19(out[19],in[19]);
	not n20(out[20],in[20]);
	not n21(out[21],in[21]);
	not n22(out[22],in[22]);
	not n23(out[23],in[23]);
	not n24(out[24],in[24]);
	not n25(out[25],in[25]);
	not n26(out[26],in[26]);
	not n27(out[27],in[27]);
	not n28(out[28],in[28]);
	not n29(out[29],in[29]);
	not n30(out[30],in[30]);
	not n31(out[31],in[31]);
	//Adder32Bit S32BAdder(out, S32Bcout, out, 32'b1);
	
endmodule

