module Mul32Bit(
	output [31:0] out,
	output cout,
	input [31:0] a,
	input [31:0] b
	);
	wire [31:0] sh0;
	wire [31:0] sh1;
	wire [31:0] sh2;
	wire [31:0] sh3;
	wire [31:0] sh4;
	wire [31:0] sh5;
	wire [31:0] sh6;
	wire [31:0] sh7;
	wire [31:0] sh8;
	wire [31:0] sh9;
	wire [31:0] sh10;
	wire [31:0] sh11;
	wire [31:0] sh12;
	wire [31:0] sh13;
	wire [31:0] sh14;
	wire [31:0] sh15;
	wire [31:0] sh16;
	wire [31:0] sh17;
	wire [31:0] sh18;
	wire [31:0] sh19;
	wire [31:0] sh20;
	wire [31:0] sh21;
	wire [31:0] sh22;
	wire [31:0] sh23;
	wire [31:0] sh24;
	wire [31:0] sh25;
	wire [31:0] sh26;
	wire [31:0] sh27;
	wire [31:0] sh28;
	wire [31:0] sh29;
	wire [31:0] sh30;
	wire [31:0] sh31;

	wire cout0;
	wire cout1;
	wire cout2;
	wire cout3;
	wire cout4;
	wire cout5;
	wire cout6;
	wire cout7;
	wire cout8;
	wire cout9;
	wire cout10;
	wire cout11;
	wire cout12;
	wire cout13;
	wire cout14;
	wire cout15;
	wire cout16;
	wire cout17;
	wire cout18;
	wire cout19;
	wire cout20;
	wire cout21;
	wire cout22;
	wire cout23;
	wire cout24;
	wire cout25;
	wire cout26;
	wire cout27;
	wire cout28;
	wire cout29;
	wire cout30;
	wire cout31;

	shiftLeft shift0(sh0,b,1'b1);
	shiftLeft shift1(sh1,sh0,1'b1);
	shiftLeft shift2(sh2,sh1,1'b1);
	shiftLeft shift3(sh3,sh2,1'b1);
	shiftLeft shift4(sh4,sh3,1'b1);
	shiftLeft shift5(sh5,sh4,1'b1);
	shiftLeft shift6(sh6,sh5,1'b1);
	shiftLeft shift7(sh7,sh6,1'b1);
	shiftLeft shift8(sh8,sh7,1'b1);
	shiftLeft shift9(sh9,sh8,1'b1);
	shiftLeft shift10(sh10,sh9,1'b1);
	shiftLeft shift11(sh11,sh10,1'b1);
	shiftLeft shift12(sh12,sh11,1'b1);
	shiftLeft shift13(sh13,sh12,1'b1);
	shiftLeft shift14(sh14,sh13,1'b1);
	shiftLeft shift15(sh15,sh14,1'b1);
	shiftLeft shift16(sh16,sh15,1'b1);
	shiftLeft shift17(sh17,sh16,1'b1);
	shiftLeft shift18(sh18,sh17,1'b1);
	shiftLeft shift19(sh19,sh18,1'b1);
	shiftLeft shift20(sh20,sh19,1'b1);
	shiftLeft shift21(sh21,sh20,1'b1);
	shiftLeft shift22(sh22,sh21,1'b1);
	shiftLeft shift23(sh23,sh22,1'b1);
	shiftLeft shift24(sh24,sh23,1'b1);
	shiftLeft shift25(sh25,sh24,1'b1);
	shiftLeft shift26(sh26,sh25,1'b1);
	shiftLeft shift27(sh27,sh26,1'b1);
	shiftLeft shift28(sh28,sh27,1'b1);
	shiftLeft shift29(sh29,sh28,1'b1);
	shiftLeft shift30(sh30,sh29,1'b1);
	shiftLeft shift31(sh31,sh30,1'b1);

and(sh0[0],sh0[0],a[0]);
and(sh0[1],sh0[1],a[0]);
and(sh0[2],sh0[2],a[0]);
and(sh0[3],sh0[3],a[0]);
and(sh0[4],sh0[4],a[0]);
and(sh0[5],sh0[5],a[0]);
and(sh0[6],sh0[6],a[0]);
and(sh0[7],sh0[7],a[0]);
and(sh0[8],sh0[8],a[0]);
and(sh0[9],sh0[9],a[0]);
and(sh0[10],sh0[10],a[0]);
and(sh0[11],sh0[11],a[0]);
and(sh0[12],sh0[12],a[0]);
and(sh0[13],sh0[13],a[0]);
and(sh0[14],sh0[14],a[0]);
and(sh0[15],sh0[15],a[0]);
and(sh0[16],sh0[16],a[0]);
and(sh0[17],sh0[17],a[0]);
and(sh0[18],sh0[18],a[0]);
and(sh0[19],sh0[19],a[0]);
and(sh0[20],sh0[20],a[0]);
and(sh0[21],sh0[21],a[0]);
and(sh0[22],sh0[22],a[0]);
and(sh0[23],sh0[23],a[0]);
and(sh0[24],sh0[24],a[0]);
and(sh0[25],sh0[25],a[0]);
and(sh0[26],sh0[26],a[0]);
and(sh0[27],sh0[27],a[0]);
and(sh0[28],sh0[28],a[0]);
and(sh0[29],sh0[29],a[0]);
and(sh0[30],sh0[30],a[0]);
and(sh0[31],sh0[31],a[0]);
and(sh1[0],sh1[0],a[1]);
and(sh1[1],sh1[1],a[1]);
and(sh1[2],sh1[2],a[1]);
and(sh1[3],sh1[3],a[1]);
and(sh1[4],sh1[4],a[1]);
and(sh1[5],sh1[5],a[1]);
and(sh1[6],sh1[6],a[1]);
and(sh1[7],sh1[7],a[1]);
and(sh1[8],sh1[8],a[1]);
and(sh1[9],sh1[9],a[1]);
and(sh1[10],sh1[10],a[1]);
and(sh1[11],sh1[11],a[1]);
and(sh1[12],sh1[12],a[1]);
and(sh1[13],sh1[13],a[1]);
and(sh1[14],sh1[14],a[1]);
and(sh1[15],sh1[15],a[1]);
and(sh1[16],sh1[16],a[1]);
and(sh1[17],sh1[17],a[1]);
and(sh1[18],sh1[18],a[1]);
and(sh1[19],sh1[19],a[1]);
and(sh1[20],sh1[20],a[1]);
and(sh1[21],sh1[21],a[1]);
and(sh1[22],sh1[22],a[1]);
and(sh1[23],sh1[23],a[1]);
and(sh1[24],sh1[24],a[1]);
and(sh1[25],sh1[25],a[1]);
and(sh1[26],sh1[26],a[1]);
and(sh1[27],sh1[27],a[1]);
and(sh1[28],sh1[28],a[1]);
and(sh1[29],sh1[29],a[1]);
and(sh1[30],sh1[30],a[1]);
and(sh1[31],sh1[31],a[1]);
and(sh2[0],sh2[0],a[2]);
and(sh2[1],sh2[1],a[2]);
and(sh2[2],sh2[2],a[2]);
and(sh2[3],sh2[3],a[2]);
and(sh2[4],sh2[4],a[2]);
and(sh2[5],sh2[5],a[2]);
and(sh2[6],sh2[6],a[2]);
and(sh2[7],sh2[7],a[2]);
and(sh2[8],sh2[8],a[2]);
and(sh2[9],sh2[9],a[2]);
and(sh2[10],sh2[10],a[2]);
and(sh2[11],sh2[11],a[2]);
and(sh2[12],sh2[12],a[2]);
and(sh2[13],sh2[13],a[2]);
and(sh2[14],sh2[14],a[2]);
and(sh2[15],sh2[15],a[2]);
and(sh2[16],sh2[16],a[2]);
and(sh2[17],sh2[17],a[2]);
and(sh2[18],sh2[18],a[2]);
and(sh2[19],sh2[19],a[2]);
and(sh2[20],sh2[20],a[2]);
and(sh2[21],sh2[21],a[2]);
and(sh2[22],sh2[22],a[2]);
and(sh2[23],sh2[23],a[2]);
and(sh2[24],sh2[24],a[2]);
and(sh2[25],sh2[25],a[2]);
and(sh2[26],sh2[26],a[2]);
and(sh2[27],sh2[27],a[2]);
and(sh2[28],sh2[28],a[2]);
and(sh2[29],sh2[29],a[2]);
and(sh2[30],sh2[30],a[2]);
and(sh2[31],sh2[31],a[2]);
and(sh3[0],sh3[0],a[3]);
and(sh3[1],sh3[1],a[3]);
and(sh3[2],sh3[2],a[3]);
and(sh3[3],sh3[3],a[3]);
and(sh3[4],sh3[4],a[3]);
and(sh3[5],sh3[5],a[3]);
and(sh3[6],sh3[6],a[3]);
and(sh3[7],sh3[7],a[3]);
and(sh3[8],sh3[8],a[3]);
and(sh3[9],sh3[9],a[3]);
and(sh3[10],sh3[10],a[3]);
and(sh3[11],sh3[11],a[3]);
and(sh3[12],sh3[12],a[3]);
and(sh3[13],sh3[13],a[3]);
and(sh3[14],sh3[14],a[3]);
and(sh3[15],sh3[15],a[3]);
and(sh3[16],sh3[16],a[3]);
and(sh3[17],sh3[17],a[3]);
and(sh3[18],sh3[18],a[3]);
and(sh3[19],sh3[19],a[3]);
and(sh3[20],sh3[20],a[3]);
and(sh3[21],sh3[21],a[3]);
and(sh3[22],sh3[22],a[3]);
and(sh3[23],sh3[23],a[3]);
and(sh3[24],sh3[24],a[3]);
and(sh3[25],sh3[25],a[3]);
and(sh3[26],sh3[26],a[3]);
and(sh3[27],sh3[27],a[3]);
and(sh3[28],sh3[28],a[3]);
and(sh3[29],sh3[29],a[3]);
and(sh3[30],sh3[30],a[3]);
and(sh3[31],sh3[31],a[3]);
and(sh4[0],sh4[0],a[4]);
and(sh4[1],sh4[1],a[4]);
and(sh4[2],sh4[2],a[4]);
and(sh4[3],sh4[3],a[4]);
and(sh4[4],sh4[4],a[4]);
and(sh4[5],sh4[5],a[4]);
and(sh4[6],sh4[6],a[4]);
and(sh4[7],sh4[7],a[4]);
and(sh4[8],sh4[8],a[4]);
and(sh4[9],sh4[9],a[4]);
and(sh4[10],sh4[10],a[4]);
and(sh4[11],sh4[11],a[4]);
and(sh4[12],sh4[12],a[4]);
and(sh4[13],sh4[13],a[4]);
and(sh4[14],sh4[14],a[4]);
and(sh4[15],sh4[15],a[4]);
and(sh4[16],sh4[16],a[4]);
and(sh4[17],sh4[17],a[4]);
and(sh4[18],sh4[18],a[4]);
and(sh4[19],sh4[19],a[4]);
and(sh4[20],sh4[20],a[4]);
and(sh4[21],sh4[21],a[4]);
and(sh4[22],sh4[22],a[4]);
and(sh4[23],sh4[23],a[4]);
and(sh4[24],sh4[24],a[4]);
and(sh4[25],sh4[25],a[4]);
and(sh4[26],sh4[26],a[4]);
and(sh4[27],sh4[27],a[4]);
and(sh4[28],sh4[28],a[4]);
and(sh4[29],sh4[29],a[4]);
and(sh4[30],sh4[30],a[4]);
and(sh4[31],sh4[31],a[4]);
and(sh5[0],sh5[0],a[5]);
and(sh5[1],sh5[1],a[5]);
and(sh5[2],sh5[2],a[5]);
and(sh5[3],sh5[3],a[5]);
and(sh5[4],sh5[4],a[5]);
and(sh5[5],sh5[5],a[5]);
and(sh5[6],sh5[6],a[5]);
and(sh5[7],sh5[7],a[5]);
and(sh5[8],sh5[8],a[5]);
and(sh5[9],sh5[9],a[5]);
and(sh5[10],sh5[10],a[5]);
and(sh5[11],sh5[11],a[5]);
and(sh5[12],sh5[12],a[5]);
and(sh5[13],sh5[13],a[5]);
and(sh5[14],sh5[14],a[5]);
and(sh5[15],sh5[15],a[5]);
and(sh5[16],sh5[16],a[5]);
and(sh5[17],sh5[17],a[5]);
and(sh5[18],sh5[18],a[5]);
and(sh5[19],sh5[19],a[5]);
and(sh5[20],sh5[20],a[5]);
and(sh5[21],sh5[21],a[5]);
and(sh5[22],sh5[22],a[5]);
and(sh5[23],sh5[23],a[5]);
and(sh5[24],sh5[24],a[5]);
and(sh5[25],sh5[25],a[5]);
and(sh5[26],sh5[26],a[5]);
and(sh5[27],sh5[27],a[5]);
and(sh5[28],sh5[28],a[5]);
and(sh5[29],sh5[29],a[5]);
and(sh5[30],sh5[30],a[5]);
and(sh5[31],sh5[31],a[5]);
and(sh6[0],sh6[0],a[6]);
and(sh6[1],sh6[1],a[6]);
and(sh6[2],sh6[2],a[6]);
and(sh6[3],sh6[3],a[6]);
and(sh6[4],sh6[4],a[6]);
and(sh6[5],sh6[5],a[6]);
and(sh6[6],sh6[6],a[6]);
and(sh6[7],sh6[7],a[6]);
and(sh6[8],sh6[8],a[6]);
and(sh6[9],sh6[9],a[6]);
and(sh6[10],sh6[10],a[6]);
and(sh6[11],sh6[11],a[6]);
and(sh6[12],sh6[12],a[6]);
and(sh6[13],sh6[13],a[6]);
and(sh6[14],sh6[14],a[6]);
and(sh6[15],sh6[15],a[6]);
and(sh6[16],sh6[16],a[6]);
and(sh6[17],sh6[17],a[6]);
and(sh6[18],sh6[18],a[6]);
and(sh6[19],sh6[19],a[6]);
and(sh6[20],sh6[20],a[6]);
and(sh6[21],sh6[21],a[6]);
and(sh6[22],sh6[22],a[6]);
and(sh6[23],sh6[23],a[6]);
and(sh6[24],sh6[24],a[6]);
and(sh6[25],sh6[25],a[6]);
and(sh6[26],sh6[26],a[6]);
and(sh6[27],sh6[27],a[6]);
and(sh6[28],sh6[28],a[6]);
and(sh6[29],sh6[29],a[6]);
and(sh6[30],sh6[30],a[6]);
and(sh6[31],sh6[31],a[6]);
and(sh7[0],sh7[0],a[7]);
and(sh7[1],sh7[1],a[7]);
and(sh7[2],sh7[2],a[7]);
and(sh7[3],sh7[3],a[7]);
and(sh7[4],sh7[4],a[7]);
and(sh7[5],sh7[5],a[7]);
and(sh7[6],sh7[6],a[7]);
and(sh7[7],sh7[7],a[7]);
and(sh7[8],sh7[8],a[7]);
and(sh7[9],sh7[9],a[7]);
and(sh7[10],sh7[10],a[7]);
and(sh7[11],sh7[11],a[7]);
and(sh7[12],sh7[12],a[7]);
and(sh7[13],sh7[13],a[7]);
and(sh7[14],sh7[14],a[7]);
and(sh7[15],sh7[15],a[7]);
and(sh7[16],sh7[16],a[7]);
and(sh7[17],sh7[17],a[7]);
and(sh7[18],sh7[18],a[7]);
and(sh7[19],sh7[19],a[7]);
and(sh7[20],sh7[20],a[7]);
and(sh7[21],sh7[21],a[7]);
and(sh7[22],sh7[22],a[7]);
and(sh7[23],sh7[23],a[7]);
and(sh7[24],sh7[24],a[7]);
and(sh7[25],sh7[25],a[7]);
and(sh7[26],sh7[26],a[7]);
and(sh7[27],sh7[27],a[7]);
and(sh7[28],sh7[28],a[7]);
and(sh7[29],sh7[29],a[7]);
and(sh7[30],sh7[30],a[7]);
and(sh7[31],sh7[31],a[7]);
and(sh8[0],sh8[0],a[8]);
and(sh8[1],sh8[1],a[8]);
and(sh8[2],sh8[2],a[8]);
and(sh8[3],sh8[3],a[8]);
and(sh8[4],sh8[4],a[8]);
and(sh8[5],sh8[5],a[8]);
and(sh8[6],sh8[6],a[8]);
and(sh8[7],sh8[7],a[8]);
and(sh8[8],sh8[8],a[8]);
and(sh8[9],sh8[9],a[8]);
and(sh8[10],sh8[10],a[8]);
and(sh8[11],sh8[11],a[8]);
and(sh8[12],sh8[12],a[8]);
and(sh8[13],sh8[13],a[8]);
and(sh8[14],sh8[14],a[8]);
and(sh8[15],sh8[15],a[8]);
and(sh8[16],sh8[16],a[8]);
and(sh8[17],sh8[17],a[8]);
and(sh8[18],sh8[18],a[8]);
and(sh8[19],sh8[19],a[8]);
and(sh8[20],sh8[20],a[8]);
and(sh8[21],sh8[21],a[8]);
and(sh8[22],sh8[22],a[8]);
and(sh8[23],sh8[23],a[8]);
and(sh8[24],sh8[24],a[8]);
and(sh8[25],sh8[25],a[8]);
and(sh8[26],sh8[26],a[8]);
and(sh8[27],sh8[27],a[8]);
and(sh8[28],sh8[28],a[8]);
and(sh8[29],sh8[29],a[8]);
and(sh8[30],sh8[30],a[8]);
and(sh8[31],sh8[31],a[8]);
and(sh9[0],sh9[0],a[9]);
and(sh9[1],sh9[1],a[9]);
and(sh9[2],sh9[2],a[9]);
and(sh9[3],sh9[3],a[9]);
and(sh9[4],sh9[4],a[9]);
and(sh9[5],sh9[5],a[9]);
and(sh9[6],sh9[6],a[9]);
and(sh9[7],sh9[7],a[9]);
and(sh9[8],sh9[8],a[9]);
and(sh9[9],sh9[9],a[9]);
and(sh9[10],sh9[10],a[9]);
and(sh9[11],sh9[11],a[9]);
and(sh9[12],sh9[12],a[9]);
and(sh9[13],sh9[13],a[9]);
and(sh9[14],sh9[14],a[9]);
and(sh9[15],sh9[15],a[9]);
and(sh9[16],sh9[16],a[9]);
and(sh9[17],sh9[17],a[9]);
and(sh9[18],sh9[18],a[9]);
and(sh9[19],sh9[19],a[9]);
and(sh9[20],sh9[20],a[9]);
and(sh9[21],sh9[21],a[9]);
and(sh9[22],sh9[22],a[9]);
and(sh9[23],sh9[23],a[9]);
and(sh9[24],sh9[24],a[9]);
and(sh9[25],sh9[25],a[9]);
and(sh9[26],sh9[26],a[9]);
and(sh9[27],sh9[27],a[9]);
and(sh9[28],sh9[28],a[9]);
and(sh9[29],sh9[29],a[9]);
and(sh9[30],sh9[30],a[9]);
and(sh9[31],sh9[31],a[9]);
and(sh10[0],sh10[0],a[10]);
and(sh10[1],sh10[1],a[10]);
and(sh10[2],sh10[2],a[10]);
and(sh10[3],sh10[3],a[10]);
and(sh10[4],sh10[4],a[10]);
and(sh10[5],sh10[5],a[10]);
and(sh10[6],sh10[6],a[10]);
and(sh10[7],sh10[7],a[10]);
and(sh10[8],sh10[8],a[10]);
and(sh10[9],sh10[9],a[10]);
and(sh10[10],sh10[10],a[10]);
and(sh10[11],sh10[11],a[10]);
and(sh10[12],sh10[12],a[10]);
and(sh10[13],sh10[13],a[10]);
and(sh10[14],sh10[14],a[10]);
and(sh10[15],sh10[15],a[10]);
and(sh10[16],sh10[16],a[10]);
and(sh10[17],sh10[17],a[10]);
and(sh10[18],sh10[18],a[10]);
and(sh10[19],sh10[19],a[10]);
and(sh10[20],sh10[20],a[10]);
and(sh10[21],sh10[21],a[10]);
and(sh10[22],sh10[22],a[10]);
and(sh10[23],sh10[23],a[10]);
and(sh10[24],sh10[24],a[10]);
and(sh10[25],sh10[25],a[10]);
and(sh10[26],sh10[26],a[10]);
and(sh10[27],sh10[27],a[10]);
and(sh10[28],sh10[28],a[10]);
and(sh10[29],sh10[29],a[10]);
and(sh10[30],sh10[30],a[10]);
and(sh10[31],sh10[31],a[10]);
and(sh11[0],sh11[0],a[11]);
and(sh11[1],sh11[1],a[11]);
and(sh11[2],sh11[2],a[11]);
and(sh11[3],sh11[3],a[11]);
and(sh11[4],sh11[4],a[11]);
and(sh11[5],sh11[5],a[11]);
and(sh11[6],sh11[6],a[11]);
and(sh11[7],sh11[7],a[11]);
and(sh11[8],sh11[8],a[11]);
and(sh11[9],sh11[9],a[11]);
and(sh11[10],sh11[10],a[11]);
and(sh11[11],sh11[11],a[11]);
and(sh11[12],sh11[12],a[11]);
and(sh11[13],sh11[13],a[11]);
and(sh11[14],sh11[14],a[11]);
and(sh11[15],sh11[15],a[11]);
and(sh11[16],sh11[16],a[11]);
and(sh11[17],sh11[17],a[11]);
and(sh11[18],sh11[18],a[11]);
and(sh11[19],sh11[19],a[11]);
and(sh11[20],sh11[20],a[11]);
and(sh11[21],sh11[21],a[11]);
and(sh11[22],sh11[22],a[11]);
and(sh11[23],sh11[23],a[11]);
and(sh11[24],sh11[24],a[11]);
and(sh11[25],sh11[25],a[11]);
and(sh11[26],sh11[26],a[11]);
and(sh11[27],sh11[27],a[11]);
and(sh11[28],sh11[28],a[11]);
and(sh11[29],sh11[29],a[11]);
and(sh11[30],sh11[30],a[11]);
and(sh11[31],sh11[31],a[11]);
and(sh12[0],sh12[0],a[12]);
and(sh12[1],sh12[1],a[12]);
and(sh12[2],sh12[2],a[12]);
and(sh12[3],sh12[3],a[12]);
and(sh12[4],sh12[4],a[12]);
and(sh12[5],sh12[5],a[12]);
and(sh12[6],sh12[6],a[12]);
and(sh12[7],sh12[7],a[12]);
and(sh12[8],sh12[8],a[12]);
and(sh12[9],sh12[9],a[12]);
and(sh12[10],sh12[10],a[12]);
and(sh12[11],sh12[11],a[12]);
and(sh12[12],sh12[12],a[12]);
and(sh12[13],sh12[13],a[12]);
and(sh12[14],sh12[14],a[12]);
and(sh12[15],sh12[15],a[12]);
and(sh12[16],sh12[16],a[12]);
and(sh12[17],sh12[17],a[12]);
and(sh12[18],sh12[18],a[12]);
and(sh12[19],sh12[19],a[12]);
and(sh12[20],sh12[20],a[12]);
and(sh12[21],sh12[21],a[12]);
and(sh12[22],sh12[22],a[12]);
and(sh12[23],sh12[23],a[12]);
and(sh12[24],sh12[24],a[12]);
and(sh12[25],sh12[25],a[12]);
and(sh12[26],sh12[26],a[12]);
and(sh12[27],sh12[27],a[12]);
and(sh12[28],sh12[28],a[12]);
and(sh12[29],sh12[29],a[12]);
and(sh12[30],sh12[30],a[12]);
and(sh12[31],sh12[31],a[12]);
and(sh13[0],sh13[0],a[13]);
and(sh13[1],sh13[1],a[13]);
and(sh13[2],sh13[2],a[13]);
and(sh13[3],sh13[3],a[13]);
and(sh13[4],sh13[4],a[13]);
and(sh13[5],sh13[5],a[13]);
and(sh13[6],sh13[6],a[13]);
and(sh13[7],sh13[7],a[13]);
and(sh13[8],sh13[8],a[13]);
and(sh13[9],sh13[9],a[13]);
and(sh13[10],sh13[10],a[13]);
and(sh13[11],sh13[11],a[13]);
and(sh13[12],sh13[12],a[13]);
and(sh13[13],sh13[13],a[13]);
and(sh13[14],sh13[14],a[13]);
and(sh13[15],sh13[15],a[13]);
and(sh13[16],sh13[16],a[13]);
and(sh13[17],sh13[17],a[13]);
and(sh13[18],sh13[18],a[13]);
and(sh13[19],sh13[19],a[13]);
and(sh13[20],sh13[20],a[13]);
and(sh13[21],sh13[21],a[13]);
and(sh13[22],sh13[22],a[13]);
and(sh13[23],sh13[23],a[13]);
and(sh13[24],sh13[24],a[13]);
and(sh13[25],sh13[25],a[13]);
and(sh13[26],sh13[26],a[13]);
and(sh13[27],sh13[27],a[13]);
and(sh13[28],sh13[28],a[13]);
and(sh13[29],sh13[29],a[13]);
and(sh13[30],sh13[30],a[13]);
and(sh13[31],sh13[31],a[13]);
and(sh14[0],sh14[0],a[14]);
and(sh14[1],sh14[1],a[14]);
and(sh14[2],sh14[2],a[14]);
and(sh14[3],sh14[3],a[14]);
and(sh14[4],sh14[4],a[14]);
and(sh14[5],sh14[5],a[14]);
and(sh14[6],sh14[6],a[14]);
and(sh14[7],sh14[7],a[14]);
and(sh14[8],sh14[8],a[14]);
and(sh14[9],sh14[9],a[14]);
and(sh14[10],sh14[10],a[14]);
and(sh14[11],sh14[11],a[14]);
and(sh14[12],sh14[12],a[14]);
and(sh14[13],sh14[13],a[14]);
and(sh14[14],sh14[14],a[14]);
and(sh14[15],sh14[15],a[14]);
and(sh14[16],sh14[16],a[14]);
and(sh14[17],sh14[17],a[14]);
and(sh14[18],sh14[18],a[14]);
and(sh14[19],sh14[19],a[14]);
and(sh14[20],sh14[20],a[14]);
and(sh14[21],sh14[21],a[14]);
and(sh14[22],sh14[22],a[14]);
and(sh14[23],sh14[23],a[14]);
and(sh14[24],sh14[24],a[14]);
and(sh14[25],sh14[25],a[14]);
and(sh14[26],sh14[26],a[14]);
and(sh14[27],sh14[27],a[14]);
and(sh14[28],sh14[28],a[14]);
and(sh14[29],sh14[29],a[14]);
and(sh14[30],sh14[30],a[14]);
and(sh14[31],sh14[31],a[14]);
and(sh15[0],sh15[0],a[15]);
and(sh15[1],sh15[1],a[15]);
and(sh15[2],sh15[2],a[15]);
and(sh15[3],sh15[3],a[15]);
and(sh15[4],sh15[4],a[15]);
and(sh15[5],sh15[5],a[15]);
and(sh15[6],sh15[6],a[15]);
and(sh15[7],sh15[7],a[15]);
and(sh15[8],sh15[8],a[15]);
and(sh15[9],sh15[9],a[15]);
and(sh15[10],sh15[10],a[15]);
and(sh15[11],sh15[11],a[15]);
and(sh15[12],sh15[12],a[15]);
and(sh15[13],sh15[13],a[15]);
and(sh15[14],sh15[14],a[15]);
and(sh15[15],sh15[15],a[15]);
and(sh15[16],sh15[16],a[15]);
and(sh15[17],sh15[17],a[15]);
and(sh15[18],sh15[18],a[15]);
and(sh15[19],sh15[19],a[15]);
and(sh15[20],sh15[20],a[15]);
and(sh15[21],sh15[21],a[15]);
and(sh15[22],sh15[22],a[15]);
and(sh15[23],sh15[23],a[15]);
and(sh15[24],sh15[24],a[15]);
and(sh15[25],sh15[25],a[15]);
and(sh15[26],sh15[26],a[15]);
and(sh15[27],sh15[27],a[15]);
and(sh15[28],sh15[28],a[15]);
and(sh15[29],sh15[29],a[15]);
and(sh15[30],sh15[30],a[15]);
and(sh15[31],sh15[31],a[15]);
and(sh16[0],sh16[0],a[16]);
and(sh16[1],sh16[1],a[16]);
and(sh16[2],sh16[2],a[16]);
and(sh16[3],sh16[3],a[16]);
and(sh16[4],sh16[4],a[16]);
and(sh16[5],sh16[5],a[16]);
and(sh16[6],sh16[6],a[16]);
and(sh16[7],sh16[7],a[16]);
and(sh16[8],sh16[8],a[16]);
and(sh16[9],sh16[9],a[16]);
and(sh16[10],sh16[10],a[16]);
and(sh16[11],sh16[11],a[16]);
and(sh16[12],sh16[12],a[16]);
and(sh16[13],sh16[13],a[16]);
and(sh16[14],sh16[14],a[16]);
and(sh16[15],sh16[15],a[16]);
and(sh16[16],sh16[16],a[16]);
and(sh16[17],sh16[17],a[16]);
and(sh16[18],sh16[18],a[16]);
and(sh16[19],sh16[19],a[16]);
and(sh16[20],sh16[20],a[16]);
and(sh16[21],sh16[21],a[16]);
and(sh16[22],sh16[22],a[16]);
and(sh16[23],sh16[23],a[16]);
and(sh16[24],sh16[24],a[16]);
and(sh16[25],sh16[25],a[16]);
and(sh16[26],sh16[26],a[16]);
and(sh16[27],sh16[27],a[16]);
and(sh16[28],sh16[28],a[16]);
and(sh16[29],sh16[29],a[16]);
and(sh16[30],sh16[30],a[16]);
and(sh16[31],sh16[31],a[16]);
and(sh17[0],sh17[0],a[17]);
and(sh17[1],sh17[1],a[17]);
and(sh17[2],sh17[2],a[17]);
and(sh17[3],sh17[3],a[17]);
and(sh17[4],sh17[4],a[17]);
and(sh17[5],sh17[5],a[17]);
and(sh17[6],sh17[6],a[17]);
and(sh17[7],sh17[7],a[17]);
and(sh17[8],sh17[8],a[17]);
and(sh17[9],sh17[9],a[17]);
and(sh17[10],sh17[10],a[17]);
and(sh17[11],sh17[11],a[17]);
and(sh17[12],sh17[12],a[17]);
and(sh17[13],sh17[13],a[17]);
and(sh17[14],sh17[14],a[17]);
and(sh17[15],sh17[15],a[17]);
and(sh17[16],sh17[16],a[17]);
and(sh17[17],sh17[17],a[17]);
and(sh17[18],sh17[18],a[17]);
and(sh17[19],sh17[19],a[17]);
and(sh17[20],sh17[20],a[17]);
and(sh17[21],sh17[21],a[17]);
and(sh17[22],sh17[22],a[17]);
and(sh17[23],sh17[23],a[17]);
and(sh17[24],sh17[24],a[17]);
and(sh17[25],sh17[25],a[17]);
and(sh17[26],sh17[26],a[17]);
and(sh17[27],sh17[27],a[17]);
and(sh17[28],sh17[28],a[17]);
and(sh17[29],sh17[29],a[17]);
and(sh17[30],sh17[30],a[17]);
and(sh17[31],sh17[31],a[17]);
and(sh18[0],sh18[0],a[18]);
and(sh18[1],sh18[1],a[18]);
and(sh18[2],sh18[2],a[18]);
and(sh18[3],sh18[3],a[18]);
and(sh18[4],sh18[4],a[18]);
and(sh18[5],sh18[5],a[18]);
and(sh18[6],sh18[6],a[18]);
and(sh18[7],sh18[7],a[18]);
and(sh18[8],sh18[8],a[18]);
and(sh18[9],sh18[9],a[18]);
and(sh18[10],sh18[10],a[18]);
and(sh18[11],sh18[11],a[18]);
and(sh18[12],sh18[12],a[18]);
and(sh18[13],sh18[13],a[18]);
and(sh18[14],sh18[14],a[18]);
and(sh18[15],sh18[15],a[18]);
and(sh18[16],sh18[16],a[18]);
and(sh18[17],sh18[17],a[18]);
and(sh18[18],sh18[18],a[18]);
and(sh18[19],sh18[19],a[18]);
and(sh18[20],sh18[20],a[18]);
and(sh18[21],sh18[21],a[18]);
and(sh18[22],sh18[22],a[18]);
and(sh18[23],sh18[23],a[18]);
and(sh18[24],sh18[24],a[18]);
and(sh18[25],sh18[25],a[18]);
and(sh18[26],sh18[26],a[18]);
and(sh18[27],sh18[27],a[18]);
and(sh18[28],sh18[28],a[18]);
and(sh18[29],sh18[29],a[18]);
and(sh18[30],sh18[30],a[18]);
and(sh18[31],sh18[31],a[18]);
and(sh19[0],sh19[0],a[19]);
and(sh19[1],sh19[1],a[19]);
and(sh19[2],sh19[2],a[19]);
and(sh19[3],sh19[3],a[19]);
and(sh19[4],sh19[4],a[19]);
and(sh19[5],sh19[5],a[19]);
and(sh19[6],sh19[6],a[19]);
and(sh19[7],sh19[7],a[19]);
and(sh19[8],sh19[8],a[19]);
and(sh19[9],sh19[9],a[19]);
and(sh19[10],sh19[10],a[19]);
and(sh19[11],sh19[11],a[19]);
and(sh19[12],sh19[12],a[19]);
and(sh19[13],sh19[13],a[19]);
and(sh19[14],sh19[14],a[19]);
and(sh19[15],sh19[15],a[19]);
and(sh19[16],sh19[16],a[19]);
and(sh19[17],sh19[17],a[19]);
and(sh19[18],sh19[18],a[19]);
and(sh19[19],sh19[19],a[19]);
and(sh19[20],sh19[20],a[19]);
and(sh19[21],sh19[21],a[19]);
and(sh19[22],sh19[22],a[19]);
and(sh19[23],sh19[23],a[19]);
and(sh19[24],sh19[24],a[19]);
and(sh19[25],sh19[25],a[19]);
and(sh19[26],sh19[26],a[19]);
and(sh19[27],sh19[27],a[19]);
and(sh19[28],sh19[28],a[19]);
and(sh19[29],sh19[29],a[19]);
and(sh19[30],sh19[30],a[19]);
and(sh19[31],sh19[31],a[19]);
and(sh20[0],sh20[0],a[20]);
and(sh20[1],sh20[1],a[20]);
and(sh20[2],sh20[2],a[20]);
and(sh20[3],sh20[3],a[20]);
and(sh20[4],sh20[4],a[20]);
and(sh20[5],sh20[5],a[20]);
and(sh20[6],sh20[6],a[20]);
and(sh20[7],sh20[7],a[20]);
and(sh20[8],sh20[8],a[20]);
and(sh20[9],sh20[9],a[20]);
and(sh20[10],sh20[10],a[20]);
and(sh20[11],sh20[11],a[20]);
and(sh20[12],sh20[12],a[20]);
and(sh20[13],sh20[13],a[20]);
and(sh20[14],sh20[14],a[20]);
and(sh20[15],sh20[15],a[20]);
and(sh20[16],sh20[16],a[20]);
and(sh20[17],sh20[17],a[20]);
and(sh20[18],sh20[18],a[20]);
and(sh20[19],sh20[19],a[20]);
and(sh20[20],sh20[20],a[20]);
and(sh20[21],sh20[21],a[20]);
and(sh20[22],sh20[22],a[20]);
and(sh20[23],sh20[23],a[20]);
and(sh20[24],sh20[24],a[20]);
and(sh20[25],sh20[25],a[20]);
and(sh20[26],sh20[26],a[20]);
and(sh20[27],sh20[27],a[20]);
and(sh20[28],sh20[28],a[20]);
and(sh20[29],sh20[29],a[20]);
and(sh20[30],sh20[30],a[20]);
and(sh20[31],sh20[31],a[20]);
and(sh21[0],sh21[0],a[21]);
and(sh21[1],sh21[1],a[21]);
and(sh21[2],sh21[2],a[21]);
and(sh21[3],sh21[3],a[21]);
and(sh21[4],sh21[4],a[21]);
and(sh21[5],sh21[5],a[21]);
and(sh21[6],sh21[6],a[21]);
and(sh21[7],sh21[7],a[21]);
and(sh21[8],sh21[8],a[21]);
and(sh21[9],sh21[9],a[21]);
and(sh21[10],sh21[10],a[21]);
and(sh21[11],sh21[11],a[21]);
and(sh21[12],sh21[12],a[21]);
and(sh21[13],sh21[13],a[21]);
and(sh21[14],sh21[14],a[21]);
and(sh21[15],sh21[15],a[21]);
and(sh21[16],sh21[16],a[21]);
and(sh21[17],sh21[17],a[21]);
and(sh21[18],sh21[18],a[21]);
and(sh21[19],sh21[19],a[21]);
and(sh21[20],sh21[20],a[21]);
and(sh21[21],sh21[21],a[21]);
and(sh21[22],sh21[22],a[21]);
and(sh21[23],sh21[23],a[21]);
and(sh21[24],sh21[24],a[21]);
and(sh21[25],sh21[25],a[21]);
and(sh21[26],sh21[26],a[21]);
and(sh21[27],sh21[27],a[21]);
and(sh21[28],sh21[28],a[21]);
and(sh21[29],sh21[29],a[21]);
and(sh21[30],sh21[30],a[21]);
and(sh21[31],sh21[31],a[21]);
and(sh22[0],sh22[0],a[22]);
and(sh22[1],sh22[1],a[22]);
and(sh22[2],sh22[2],a[22]);
and(sh22[3],sh22[3],a[22]);
and(sh22[4],sh22[4],a[22]);
and(sh22[5],sh22[5],a[22]);
and(sh22[6],sh22[6],a[22]);
and(sh22[7],sh22[7],a[22]);
and(sh22[8],sh22[8],a[22]);
and(sh22[9],sh22[9],a[22]);
and(sh22[10],sh22[10],a[22]);
and(sh22[11],sh22[11],a[22]);
and(sh22[12],sh22[12],a[22]);
and(sh22[13],sh22[13],a[22]);
and(sh22[14],sh22[14],a[22]);
and(sh22[15],sh22[15],a[22]);
and(sh22[16],sh22[16],a[22]);
and(sh22[17],sh22[17],a[22]);
and(sh22[18],sh22[18],a[22]);
and(sh22[19],sh22[19],a[22]);
and(sh22[20],sh22[20],a[22]);
and(sh22[21],sh22[21],a[22]);
and(sh22[22],sh22[22],a[22]);
and(sh22[23],sh22[23],a[22]);
and(sh22[24],sh22[24],a[22]);
and(sh22[25],sh22[25],a[22]);
and(sh22[26],sh22[26],a[22]);
and(sh22[27],sh22[27],a[22]);
and(sh22[28],sh22[28],a[22]);
and(sh22[29],sh22[29],a[22]);
and(sh22[30],sh22[30],a[22]);
and(sh22[31],sh22[31],a[22]);
and(sh23[0],sh23[0],a[23]);
and(sh23[1],sh23[1],a[23]);
and(sh23[2],sh23[2],a[23]);
and(sh23[3],sh23[3],a[23]);
and(sh23[4],sh23[4],a[23]);
and(sh23[5],sh23[5],a[23]);
and(sh23[6],sh23[6],a[23]);
and(sh23[7],sh23[7],a[23]);
and(sh23[8],sh23[8],a[23]);
and(sh23[9],sh23[9],a[23]);
and(sh23[10],sh23[10],a[23]);
and(sh23[11],sh23[11],a[23]);
and(sh23[12],sh23[12],a[23]);
and(sh23[13],sh23[13],a[23]);
and(sh23[14],sh23[14],a[23]);
and(sh23[15],sh23[15],a[23]);
and(sh23[16],sh23[16],a[23]);
and(sh23[17],sh23[17],a[23]);
and(sh23[18],sh23[18],a[23]);
and(sh23[19],sh23[19],a[23]);
and(sh23[20],sh23[20],a[23]);
and(sh23[21],sh23[21],a[23]);
and(sh23[22],sh23[22],a[23]);
and(sh23[23],sh23[23],a[23]);
and(sh23[24],sh23[24],a[23]);
and(sh23[25],sh23[25],a[23]);
and(sh23[26],sh23[26],a[23]);
and(sh23[27],sh23[27],a[23]);
and(sh23[28],sh23[28],a[23]);
and(sh23[29],sh23[29],a[23]);
and(sh23[30],sh23[30],a[23]);
and(sh23[31],sh23[31],a[23]);
and(sh24[0],sh24[0],a[24]);
and(sh24[1],sh24[1],a[24]);
and(sh24[2],sh24[2],a[24]);
and(sh24[3],sh24[3],a[24]);
and(sh24[4],sh24[4],a[24]);
and(sh24[5],sh24[5],a[24]);
and(sh24[6],sh24[6],a[24]);
and(sh24[7],sh24[7],a[24]);
and(sh24[8],sh24[8],a[24]);
and(sh24[9],sh24[9],a[24]);
and(sh24[10],sh24[10],a[24]);
and(sh24[11],sh24[11],a[24]);
and(sh24[12],sh24[12],a[24]);
and(sh24[13],sh24[13],a[24]);
and(sh24[14],sh24[14],a[24]);
and(sh24[15],sh24[15],a[24]);
and(sh24[16],sh24[16],a[24]);
and(sh24[17],sh24[17],a[24]);
and(sh24[18],sh24[18],a[24]);
and(sh24[19],sh24[19],a[24]);
and(sh24[20],sh24[20],a[24]);
and(sh24[21],sh24[21],a[24]);
and(sh24[22],sh24[22],a[24]);
and(sh24[23],sh24[23],a[24]);
and(sh24[24],sh24[24],a[24]);
and(sh24[25],sh24[25],a[24]);
and(sh24[26],sh24[26],a[24]);
and(sh24[27],sh24[27],a[24]);
and(sh24[28],sh24[28],a[24]);
and(sh24[29],sh24[29],a[24]);
and(sh24[30],sh24[30],a[24]);
and(sh24[31],sh24[31],a[24]);
and(sh25[0],sh25[0],a[25]);
and(sh25[1],sh25[1],a[25]);
and(sh25[2],sh25[2],a[25]);
and(sh25[3],sh25[3],a[25]);
and(sh25[4],sh25[4],a[25]);
and(sh25[5],sh25[5],a[25]);
and(sh25[6],sh25[6],a[25]);
and(sh25[7],sh25[7],a[25]);
and(sh25[8],sh25[8],a[25]);
and(sh25[9],sh25[9],a[25]);
and(sh25[10],sh25[10],a[25]);
and(sh25[11],sh25[11],a[25]);
and(sh25[12],sh25[12],a[25]);
and(sh25[13],sh25[13],a[25]);
and(sh25[14],sh25[14],a[25]);
and(sh25[15],sh25[15],a[25]);
and(sh25[16],sh25[16],a[25]);
and(sh25[17],sh25[17],a[25]);
and(sh25[18],sh25[18],a[25]);
and(sh25[19],sh25[19],a[25]);
and(sh25[20],sh25[20],a[25]);
and(sh25[21],sh25[21],a[25]);
and(sh25[22],sh25[22],a[25]);
and(sh25[23],sh25[23],a[25]);
and(sh25[24],sh25[24],a[25]);
and(sh25[25],sh25[25],a[25]);
and(sh25[26],sh25[26],a[25]);
and(sh25[27],sh25[27],a[25]);
and(sh25[28],sh25[28],a[25]);
and(sh25[29],sh25[29],a[25]);
and(sh25[30],sh25[30],a[25]);
and(sh25[31],sh25[31],a[25]);
and(sh26[0],sh26[0],a[26]);
and(sh26[1],sh26[1],a[26]);
and(sh26[2],sh26[2],a[26]);
and(sh26[3],sh26[3],a[26]);
and(sh26[4],sh26[4],a[26]);
and(sh26[5],sh26[5],a[26]);
and(sh26[6],sh26[6],a[26]);
and(sh26[7],sh26[7],a[26]);
and(sh26[8],sh26[8],a[26]);
and(sh26[9],sh26[9],a[26]);
and(sh26[10],sh26[10],a[26]);
and(sh26[11],sh26[11],a[26]);
and(sh26[12],sh26[12],a[26]);
and(sh26[13],sh26[13],a[26]);
and(sh26[14],sh26[14],a[26]);
and(sh26[15],sh26[15],a[26]);
and(sh26[16],sh26[16],a[26]);
and(sh26[17],sh26[17],a[26]);
and(sh26[18],sh26[18],a[26]);
and(sh26[19],sh26[19],a[26]);
and(sh26[20],sh26[20],a[26]);
and(sh26[21],sh26[21],a[26]);
and(sh26[22],sh26[22],a[26]);
and(sh26[23],sh26[23],a[26]);
and(sh26[24],sh26[24],a[26]);
and(sh26[25],sh26[25],a[26]);
and(sh26[26],sh26[26],a[26]);
and(sh26[27],sh26[27],a[26]);
and(sh26[28],sh26[28],a[26]);
and(sh26[29],sh26[29],a[26]);
and(sh26[30],sh26[30],a[26]);
and(sh26[31],sh26[31],a[26]);
and(sh27[0],sh27[0],a[27]);
and(sh27[1],sh27[1],a[27]);
and(sh27[2],sh27[2],a[27]);
and(sh27[3],sh27[3],a[27]);
and(sh27[4],sh27[4],a[27]);
and(sh27[5],sh27[5],a[27]);
and(sh27[6],sh27[6],a[27]);
and(sh27[7],sh27[7],a[27]);
and(sh27[8],sh27[8],a[27]);
and(sh27[9],sh27[9],a[27]);
and(sh27[10],sh27[10],a[27]);
and(sh27[11],sh27[11],a[27]);
and(sh27[12],sh27[12],a[27]);
and(sh27[13],sh27[13],a[27]);
and(sh27[14],sh27[14],a[27]);
and(sh27[15],sh27[15],a[27]);
and(sh27[16],sh27[16],a[27]);
and(sh27[17],sh27[17],a[27]);
and(sh27[18],sh27[18],a[27]);
and(sh27[19],sh27[19],a[27]);
and(sh27[20],sh27[20],a[27]);
and(sh27[21],sh27[21],a[27]);
and(sh27[22],sh27[22],a[27]);
and(sh27[23],sh27[23],a[27]);
and(sh27[24],sh27[24],a[27]);
and(sh27[25],sh27[25],a[27]);
and(sh27[26],sh27[26],a[27]);
and(sh27[27],sh27[27],a[27]);
and(sh27[28],sh27[28],a[27]);
and(sh27[29],sh27[29],a[27]);
and(sh27[30],sh27[30],a[27]);
and(sh27[31],sh27[31],a[27]);
and(sh28[0],sh28[0],a[28]);
and(sh28[1],sh28[1],a[28]);
and(sh28[2],sh28[2],a[28]);
and(sh28[3],sh28[3],a[28]);
and(sh28[4],sh28[4],a[28]);
and(sh28[5],sh28[5],a[28]);
and(sh28[6],sh28[6],a[28]);
and(sh28[7],sh28[7],a[28]);
and(sh28[8],sh28[8],a[28]);
and(sh28[9],sh28[9],a[28]);
and(sh28[10],sh28[10],a[28]);
and(sh28[11],sh28[11],a[28]);
and(sh28[12],sh28[12],a[28]);
and(sh28[13],sh28[13],a[28]);
and(sh28[14],sh28[14],a[28]);
and(sh28[15],sh28[15],a[28]);
and(sh28[16],sh28[16],a[28]);
and(sh28[17],sh28[17],a[28]);
and(sh28[18],sh28[18],a[28]);
and(sh28[19],sh28[19],a[28]);
and(sh28[20],sh28[20],a[28]);
and(sh28[21],sh28[21],a[28]);
and(sh28[22],sh28[22],a[28]);
and(sh28[23],sh28[23],a[28]);
and(sh28[24],sh28[24],a[28]);
and(sh28[25],sh28[25],a[28]);
and(sh28[26],sh28[26],a[28]);
and(sh28[27],sh28[27],a[28]);
and(sh28[28],sh28[28],a[28]);
and(sh28[29],sh28[29],a[28]);
and(sh28[30],sh28[30],a[28]);
and(sh28[31],sh28[31],a[28]);
and(sh29[0],sh29[0],a[29]);
and(sh29[1],sh29[1],a[29]);
and(sh29[2],sh29[2],a[29]);
and(sh29[3],sh29[3],a[29]);
and(sh29[4],sh29[4],a[29]);
and(sh29[5],sh29[5],a[29]);
and(sh29[6],sh29[6],a[29]);
and(sh29[7],sh29[7],a[29]);
and(sh29[8],sh29[8],a[29]);
and(sh29[9],sh29[9],a[29]);
and(sh29[10],sh29[10],a[29]);
and(sh29[11],sh29[11],a[29]);
and(sh29[12],sh29[12],a[29]);
and(sh29[13],sh29[13],a[29]);
and(sh29[14],sh29[14],a[29]);
and(sh29[15],sh29[15],a[29]);
and(sh29[16],sh29[16],a[29]);
and(sh29[17],sh29[17],a[29]);
and(sh29[18],sh29[18],a[29]);
and(sh29[19],sh29[19],a[29]);
and(sh29[20],sh29[20],a[29]);
and(sh29[21],sh29[21],a[29]);
and(sh29[22],sh29[22],a[29]);
and(sh29[23],sh29[23],a[29]);
and(sh29[24],sh29[24],a[29]);
and(sh29[25],sh29[25],a[29]);
and(sh29[26],sh29[26],a[29]);
and(sh29[27],sh29[27],a[29]);
and(sh29[28],sh29[28],a[29]);
and(sh29[29],sh29[29],a[29]);
and(sh29[30],sh29[30],a[29]);
and(sh29[31],sh29[31],a[29]);
and(sh30[0],sh30[0],a[30]);
and(sh30[1],sh30[1],a[30]);
and(sh30[2],sh30[2],a[30]);
and(sh30[3],sh30[3],a[30]);
and(sh30[4],sh30[4],a[30]);
and(sh30[5],sh30[5],a[30]);
and(sh30[6],sh30[6],a[30]);
and(sh30[7],sh30[7],a[30]);
and(sh30[8],sh30[8],a[30]);
and(sh30[9],sh30[9],a[30]);
and(sh30[10],sh30[10],a[30]);
and(sh30[11],sh30[11],a[30]);
and(sh30[12],sh30[12],a[30]);
and(sh30[13],sh30[13],a[30]);
and(sh30[14],sh30[14],a[30]);
and(sh30[15],sh30[15],a[30]);
and(sh30[16],sh30[16],a[30]);
and(sh30[17],sh30[17],a[30]);
and(sh30[18],sh30[18],a[30]);
and(sh30[19],sh30[19],a[30]);
and(sh30[20],sh30[20],a[30]);
and(sh30[21],sh30[21],a[30]);
and(sh30[22],sh30[22],a[30]);
and(sh30[23],sh30[23],a[30]);
and(sh30[24],sh30[24],a[30]);
and(sh30[25],sh30[25],a[30]);
and(sh30[26],sh30[26],a[30]);
and(sh30[27],sh30[27],a[30]);
and(sh30[28],sh30[28],a[30]);
and(sh30[29],sh30[29],a[30]);
and(sh30[30],sh30[30],a[30]);
and(sh30[31],sh30[31],a[30]);
and(sh31[0],sh31[0],a[31]);
and(sh31[1],sh31[1],a[31]);
and(sh31[2],sh31[2],a[31]);
and(sh31[3],sh31[3],a[31]);
and(sh31[4],sh31[4],a[31]);
and(sh31[5],sh31[5],a[31]);
and(sh31[6],sh31[6],a[31]);
and(sh31[7],sh31[7],a[31]);
and(sh31[8],sh31[8],a[31]);
and(sh31[9],sh31[9],a[31]);
and(sh31[10],sh31[10],a[31]);
and(sh31[11],sh31[11],a[31]);
and(sh31[12],sh31[12],a[31]);
and(sh31[13],sh31[13],a[31]);
and(sh31[14],sh31[14],a[31]);
and(sh31[15],sh31[15],a[31]);
and(sh31[16],sh31[16],a[31]);
and(sh31[17],sh31[17],a[31]);
and(sh31[18],sh31[18],a[31]);
and(sh31[19],sh31[19],a[31]);
and(sh31[20],sh31[20],a[31]);
and(sh31[21],sh31[21],a[31]);
and(sh31[22],sh31[22],a[31]);
and(sh31[23],sh31[23],a[31]);
and(sh31[24],sh31[24],a[31]);
and(sh31[25],sh31[25],a[31]);
and(sh31[26],sh31[26],a[31]);
and(sh31[27],sh31[27],a[31]);
and(sh31[28],sh31[28],a[31]);
and(sh31[29],sh31[29],a[31]);
and(sh31[30],sh31[30],a[31]);
and(sh31[31],sh31[31],a[31]);


	Adder32Bit add0(out,cout0,sh1,sh0);
	Adder32Bit add1(out,cout1,out,sh1);
	Adder32Bit add2(out,cout2,out,sh2);
	Adder32Bit add3(out,cout3,out,sh3);
	Adder32Bit add4(out,cout4,out,sh4);
	Adder32Bit add5(out,cout5,out,sh5);
	Adder32Bit add6(out,cout6,out,sh6);
	Adder32Bit add7(out,cout7,out,sh7);
	Adder32Bit add8(out,cout8,out,sh8);
	Adder32Bit add9(out,cout9,out,sh9);
	Adder32Bit add10(out,cout10,out,sh10);
	Adder32Bit add11(out,cout11,out,sh11);
	Adder32Bit add12(out,cout12,out,sh12);
	Adder32Bit add13(out,cout13,out,sh13);
	Adder32Bit add14(out,cout14,out,sh14);
	Adder32Bit add15(out,cout15,out,sh15);
	Adder32Bit add16(out,cout16,out,sh16);
	Adder32Bit add17(out,cout17,out,sh17);
	Adder32Bit add18(out,cout18,out,sh18);
	Adder32Bit add19(out,cout19,out,sh19);
	Adder32Bit add20(out,cout20,out,sh20);
	Adder32Bit add21(out,cout21,out,sh21);
	Adder32Bit add22(out,cout22,out,sh22);
	Adder32Bit add23(out,cout23,out,sh23);
	Adder32Bit add24(out,cout24,out,sh24);
	Adder32Bit add25(out,cout25,out,sh25);
	Adder32Bit add26(out,cout26,out,sh26);
	Adder32Bit add27(out,cout27,out,sh27);
	Adder32Bit add28(out,cout28,out,sh28);
	Adder32Bit add29(out,cout29,out,sh29);
	Adder32Bit add30(out,cout30,out,sh30);
	Adder32Bit add31(out,cout31,out,sh31);

	//or(cout,cout0,cout1,cout2,cout3,cout4,cout5,cout6,cout7,cout8,cout9,cout10,cout11,cout12,cout13,cout14,cout15,cout16,cout17,cout18,cout19,cout20,cout21,cout22,cout23,cout24,cout25,cout26,cout27,cout28,cout29,cout30,cout31);

endmodule
